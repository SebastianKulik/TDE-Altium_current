*****************************************************************************
** LM5116_BUCK_BLOCK.WB_LM5116_BUCK_BLOCK_WITH_RRAMP.D1 Spice Model
*****************************************************************************
** (C) Copyright 2016 Texas Instruments Incorporated. All rights reserved.
** This model is designed as an aid for customers of Texas Instruments.
** TI and its licensors and suppliers make no warranties, either expressed
** or implied, with respect to this model, including the warranties of
** merchantability or fitness for a particular purpose. The model is
** provided solely on an "as is" basis. The entire risk as to its quality
** and performance is with the customer
*****************************************************************************
*****************************************************************************

.subckt LM5116_BUCK_BLOCK_WB_LM5116_BUCK_BLOCK_WITH_RRAMP_D1_ENCR 10 11
.include isspice://../LM5116_BUCK_BLOCK.WB_LM5116_BUCK_BLOCK_WITH_RRAMP.D1.enl
XCALL 10 11 LM5116_BUCK_BLOCK_WB_LM5116_BUCK_BLOCK_WITH_RRAMP_D1 
.ENDS
