***********************************
*     Created by WB Importer      *
***********************************
.subckt LM5116_BUCK_BLOCK_WB_LM5116_BUCK_BLOCK_WITH_RRAMP_Cvcc 10 0
Cvcc 10 0 1.0E-6

.ends
