***********************************
*     Created by WB Importer      *
***********************************
.subckt LM5116_BUCK_BLOCK_WB_LM5116_BUCK_BLOCK_WITH_RRAMP_Ccomp 8 24
Ccomp 8 24 1.0E-9

.ends
