***********************************
*     Created by WB Importer      *
***********************************
.SUBCKT LM5116_BUCK_BLOCK_Cout_WB_CAP_AL 2 4
R1 2 3 0.44
C1 3 1 2.7E-5 IC = 0.0
R3 5 4 150; free space reduced by sqrt(dielectric constant)
R2 2 4 3.703703703703704E7
R4 3 26 5.5E10
R6 3 7 55000.0
C5 7 1 1.08E-5 IC = 0.0
R7 3 10 55000.0
C6 10 1 1.08E-5 IC = 0.0
R8 3 13 55000.0
C7 13 1 1.08E-5 IC = 0.0
C2 26 1 1.08E-5 IC = 0.0
R9 3 28 5.5E8
C3 28 1 1.08E-5 IC = 0.0
R10 3 29 5500000.0
C4 29 1 1.08E-5 IC = 0.0
L8 1 5 0.2e-9
R24 1 5 1.32
L12 5 4 10e-12
.ENDS
