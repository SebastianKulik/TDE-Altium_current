***********************************
*     Created by WB Importer      *
***********************************
.subckt LM5116_BUCK_BLOCK_WB_LM5116_BUCK_BLOCK_WITH_RRAMP_Rsense 12 0
Rsense 12 0 0.025

.ends
