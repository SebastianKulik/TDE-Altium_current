*****************************************************************************
** LM5116_BUCK_BLOCK.U1.WB_LM5116 Spice Model
*****************************************************************************
** (C) Copyright 2016 Texas Instruments Incorporated. All rights reserved.
** This model is designed as an aid for customers of Texas Instruments.
** TI and its licensors and suppliers make no warranties, either expressed
** or implied, with respect to this model, including the warranties of
** merchantability or fitness for a particular purpose. The model is
** provided solely on an "as is" basis. The entire risk as to its quality
** and performance is with the customer
*****************************************************************************
*****************************************************************************

.SUBCKT LM5116_BUCK_BLOCK_U1_WB_LM5116_ENCR VIN UVLO RT EN RAMP GND SS FB COMP OUT DEMB CS CSG PGND LO VCC VCCX BST HO SW
.include isspice://../LM5116_BUCK_BLOCK.U1.WB_LM5116.enl
XCALL VIN UVLO RT EN RAMP GND SS FB COMP OUT DEMB CS CSG PGND LO VCC VCCX BST HO SW LM5116_BUCK_BLOCK_U1_WB_LM5116 
.ENDS
