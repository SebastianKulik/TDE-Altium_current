***********************************
*     Created by WB Importer      *
***********************************
.subckt LM5116_BUCK_BLOCK_WB_LM5116_BUCK_BLOCK_WITH_RRAMP_Ruv1 2 0
Ruv1 2 0 3400.0

.ends
