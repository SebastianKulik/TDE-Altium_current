***********************************
*     Created by WB Importer      *
***********************************
.SUBCKT LM5116_BUCK_BLOCK_L1_WB_INDUCTOR 1 2
*{ L = 1.0E-4 DCR = 0.106 }
* PARAMETERS: L INDUCTANCE IN HENRIES, DCR DC SERIES RESISTANCE IN OHMS

L1 2 3 1.0E-4
RDCR 3 1 0.106

.ENDS
